module ip2;
  ip4 u_ip4 ();
endmodule
