module ip1;
endmodule
