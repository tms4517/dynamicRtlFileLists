module ip4;
endmodule
