module ip3;
endmodule
