module ip2;
endmodule
