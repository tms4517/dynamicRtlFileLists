module ip1;
  ip3 u_ip3 ();
endmodule
