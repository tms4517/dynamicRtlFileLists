module top;
    ip1 u_ip1 ();
    ip2 u_ip2 ();
endmodule
